magic
tech sky130A
timestamp 1701680991
<< error_p >>
rect -60 -20 110 120
<< nwell >>
rect -60 -20 110 120
<< pmos >>
rect 0 0 50 100
<< pdiff >>
rect -40 90 0 100
rect -40 70 -30 90
rect -10 70 0 90
rect -40 30 0 70
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 90 90 100
rect 50 70 60 90
rect 80 70 90 90
rect 50 30 90 70
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
<< pdiffc >>
rect -30 70 -10 90
rect -30 10 -10 30
rect 60 70 80 90
rect 60 10 80 30
<< poly >>
rect 0 100 50 115
rect 0 -15 50 0
<< locali >>
rect -40 90 0 100
rect -40 70 -30 90
rect -10 70 0 90
rect -40 30 0 70
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 50 90 90 100
rect 50 70 60 90
rect 80 70 90 90
rect 50 30 90 70
rect 50 10 60 30
rect 80 10 90 30
rect 50 0 90 10
<< end >>
