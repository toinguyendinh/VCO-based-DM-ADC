magic
tech sky130A
timestamp 1701680991
<< error_p >>
rect -40 0 0 200
rect 130 0 170 200
<< nmos >>
rect 0 0 130 200
<< ndiff >>
rect -40 190 0 200
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 130 190 170 200
rect 130 170 140 190
rect 160 170 170 190
rect 130 150 170 170
rect 130 130 140 150
rect 160 130 170 150
rect 130 110 170 130
rect 130 90 140 110
rect 160 90 170 110
rect 130 70 170 90
rect 130 50 140 70
rect 160 50 170 70
rect 130 30 170 50
rect 130 10 140 30
rect 160 10 170 30
rect 130 0 170 10
<< ndiffc >>
rect -30 170 -10 190
rect -30 130 -10 150
rect -30 90 -10 110
rect -30 50 -10 70
rect -30 10 -10 30
rect 140 170 160 190
rect 140 130 160 150
rect 140 90 160 110
rect 140 50 160 70
rect 140 10 160 30
<< poly >>
rect 0 200 130 220
rect 0 -20 130 0
<< locali >>
rect -40 190 0 200
rect -40 170 -30 190
rect -10 170 0 190
rect -40 150 0 170
rect -40 130 -30 150
rect -10 130 0 150
rect -40 110 0 130
rect -40 90 -30 110
rect -10 90 0 110
rect -40 70 0 90
rect -40 50 -30 70
rect -10 50 0 70
rect -40 30 0 50
rect -40 10 -30 30
rect -10 10 0 30
rect -40 0 0 10
rect 130 190 170 200
rect 130 170 140 190
rect 160 170 170 190
rect 130 150 170 170
rect 130 130 140 150
rect 160 130 170 150
rect 130 110 170 130
rect 130 90 140 110
rect 160 90 170 110
rect 130 70 170 90
rect 130 50 140 70
rect 160 50 170 70
rect 130 30 170 50
rect 130 10 140 30
rect 160 10 170 30
rect 130 0 170 10
<< end >>
