magic
tech sky130A
timestamp 1701680991
<< error_p >>
rect -60 220 190 680
<< nwell >>
rect -60 220 190 680
<< pmos >>
rect 0 250 130 650
<< pdiff >>
rect -40 640 0 650
rect -40 620 -30 640
rect -10 620 0 640
rect -40 600 0 620
rect -40 580 -30 600
rect -10 580 0 600
rect -40 560 0 580
rect -40 540 -30 560
rect -10 540 0 560
rect -40 520 0 540
rect -40 500 -30 520
rect -10 500 0 520
rect -40 480 0 500
rect -40 460 -30 480
rect -10 460 0 480
rect -40 440 0 460
rect -40 420 -30 440
rect -10 420 0 440
rect -40 400 0 420
rect -40 380 -30 400
rect -10 380 0 400
rect -40 360 0 380
rect -40 340 -30 360
rect -10 340 0 360
rect -40 320 0 340
rect -40 300 -30 320
rect -10 300 0 320
rect -40 280 0 300
rect -40 260 -30 280
rect -10 260 0 280
rect -40 250 0 260
rect 130 640 170 650
rect 130 620 140 640
rect 160 620 170 640
rect 130 600 170 620
rect 130 580 140 600
rect 160 580 170 600
rect 130 560 170 580
rect 130 540 140 560
rect 160 540 170 560
rect 130 520 170 540
rect 130 500 140 520
rect 160 500 170 520
rect 130 480 170 500
rect 130 460 140 480
rect 160 460 170 480
rect 130 440 170 460
rect 130 420 140 440
rect 160 420 170 440
rect 130 400 170 420
rect 130 380 140 400
rect 160 380 170 400
rect 130 360 170 380
rect 130 340 140 360
rect 160 340 170 360
rect 130 320 170 340
rect 130 300 140 320
rect 160 300 170 320
rect 130 280 170 300
rect 130 260 140 280
rect 160 260 170 280
rect 130 250 170 260
<< pdiffc >>
rect -30 620 -10 640
rect -30 580 -10 600
rect -30 540 -10 560
rect -30 500 -10 520
rect -30 460 -10 480
rect -30 420 -10 440
rect -30 380 -10 400
rect -30 340 -10 360
rect -30 300 -10 320
rect -30 260 -10 280
rect 140 620 160 640
rect 140 580 160 600
rect 140 540 160 560
rect 140 500 160 520
rect 140 460 160 480
rect 140 420 160 440
rect 140 380 160 400
rect 140 340 160 360
rect 140 300 160 320
rect 140 260 160 280
<< poly >>
rect 0 650 130 670
rect 0 230 130 250
<< locali >>
rect -40 640 0 650
rect -40 620 -30 640
rect -10 620 0 640
rect -40 600 0 620
rect -40 580 -30 600
rect -10 580 0 600
rect -40 560 0 580
rect -40 540 -30 560
rect -10 540 0 560
rect -40 520 0 540
rect -40 500 -30 520
rect -10 500 0 520
rect -40 480 0 500
rect -40 460 -30 480
rect -10 460 0 480
rect -40 440 0 460
rect -40 420 -30 440
rect -10 420 0 440
rect -40 400 0 420
rect -40 380 -30 400
rect -10 380 0 400
rect -40 360 0 380
rect -40 340 -30 360
rect -10 340 0 360
rect -40 320 0 340
rect -40 300 -30 320
rect -10 300 0 320
rect -40 280 0 300
rect -40 260 -30 280
rect -10 260 0 280
rect -40 250 0 260
rect 130 640 170 650
rect 130 620 140 640
rect 160 620 170 640
rect 130 600 170 620
rect 130 580 140 600
rect 160 580 170 600
rect 130 560 170 580
rect 130 540 140 560
rect 160 540 170 560
rect 130 520 170 540
rect 130 500 140 520
rect 160 500 170 520
rect 130 480 170 500
rect 130 460 140 480
rect 160 460 170 480
rect 130 440 170 460
rect 130 420 140 440
rect 160 420 170 440
rect 130 400 170 420
rect 130 380 140 400
rect 160 380 170 400
rect 130 360 170 380
rect 130 340 140 360
rect 160 340 170 360
rect 130 320 170 340
rect 130 300 140 320
rect 160 300 170 320
rect 130 280 170 300
rect 130 260 140 280
rect 160 260 170 280
rect 130 250 170 260
<< end >>
